module xbar_sys_1_15 #(
        // parameter NM = 1,
        // parameter NS = 16
    )(
    (* X_INTERFACE_PARAMETER = "XIL_INTERFACENAME s_axi_clk, ASSOCIATED_BUSIF s_axi_0:m_axi_0:m_axi_1:m_axi_2:m_axi_3:m_axi_4:m_axi_5:m_axi_6:m_axi_7:m_axi_8:m_axi_9:m_axi_10:m_axi_11:m_axi_12:m_axi_13:m_axi_14:m_axi_15, ASSOCIATED_RESET s_axi_aresetn" *)
    (* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 s_axi_clk CLK" *)
    input wire S_AXI_ACLK,
    (* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 s_axi_aresetn RST" *)
    input wire S_AXI_ARESETN,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 AWVALID" *)
    output wire M_AXI_0_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 AWREADY" *)
    input wire M_AXI_0_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 AWADDR" *)
    output wire [32-1:0] M_AXI_0_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 AWPROT" *)
    output wire [2:0] M_AXI_0_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 WVALID" *)
    output wire M_AXI_0_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 WREADY" *)
    input wire M_AXI_0_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 WDATA" *)
    output wire [32-1:0] M_AXI_0_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 WSTRB" *)
    output wire [4-1:0] M_AXI_0_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 BVALID" *)
    input wire M_AXI_0_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 BREADY" *)
    output wire M_AXI_0_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 BRESP" *)
    input wire [1:0] M_AXI_0_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 ARVALID" *)
    output wire M_AXI_0_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 ARREADY" *)
    input wire M_AXI_0_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 ARADDR" *)
    output wire [32-1:0] M_AXI_0_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 ARPROT" *)
    output wire [2:0] M_AXI_0_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 RVALID" *)
    input wire M_AXI_0_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 RREADY" *)
    output wire M_AXI_0_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 RRESP" *)
    input wire [1:0] M_AXI_0_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_0 RDATA" *)
    input wire [32-1:0] M_AXI_0_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 AWVALID" *)
    output wire M_AXI_1_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 AWREADY" *)
    input wire M_AXI_1_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 AWADDR" *)
    output wire [32-1:0] M_AXI_1_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 AWPROT" *)
    output wire [2:0] M_AXI_1_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 WVALID" *)
    output wire M_AXI_1_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 WREADY" *)
    input wire M_AXI_1_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 WDATA" *)
    output wire [32-1:0] M_AXI_1_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 WSTRB" *)
    output wire [4-1:0] M_AXI_1_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 BVALID" *)
    input wire M_AXI_1_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 BREADY" *)
    output wire M_AXI_1_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 BRESP" *)
    input wire [1:0] M_AXI_1_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 ARVALID" *)
    output wire M_AXI_1_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 ARREADY" *)
    input wire M_AXI_1_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 ARADDR" *)
    output wire [32-1:0] M_AXI_1_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 ARPROT" *)
    output wire [2:0] M_AXI_1_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 RVALID" *)
    input wire M_AXI_1_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 RREADY" *)
    output wire M_AXI_1_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 RRESP" *)
    input wire [1:0] M_AXI_1_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_1 RDATA" *)
    input wire [32-1:0] M_AXI_1_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 AWVALID" *)
    output wire M_AXI_2_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 AWREADY" *)
    input wire M_AXI_2_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 AWADDR" *)
    output wire [32-1:0] M_AXI_2_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 AWPROT" *)
    output wire [2:0] M_AXI_2_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 WVALID" *)
    output wire M_AXI_2_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 WREADY" *)
    input wire M_AXI_2_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 WDATA" *)
    output wire [32-1:0] M_AXI_2_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 WSTRB" *)
    output wire [4-1:0] M_AXI_2_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 BVALID" *)
    input wire M_AXI_2_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 BREADY" *)
    output wire M_AXI_2_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 BRESP" *)
    input wire [1:0] M_AXI_2_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 ARVALID" *)
    output wire M_AXI_2_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 ARREADY" *)
    input wire M_AXI_2_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 ARADDR" *)
    output wire [32-1:0] M_AXI_2_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 ARPROT" *)
    output wire [2:0] M_AXI_2_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 RVALID" *)
    input wire M_AXI_2_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 RREADY" *)
    output wire M_AXI_2_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 RRESP" *)
    input wire [1:0] M_AXI_2_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_2 RDATA" *)
    input wire [32-1:0] M_AXI_2_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 AWVALID" *)
    output wire M_AXI_3_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 AWREADY" *)
    input wire M_AXI_3_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 AWADDR" *)
    output wire [32-1:0] M_AXI_3_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 AWPROT" *)
    output wire [2:0] M_AXI_3_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 WVALID" *)
    output wire M_AXI_3_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 WREADY" *)
    input wire M_AXI_3_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 WDATA" *)
    output wire [32-1:0] M_AXI_3_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 WSTRB" *)
    output wire [4-1:0] M_AXI_3_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 BVALID" *)
    input wire M_AXI_3_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 BREADY" *)
    output wire M_AXI_3_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 BRESP" *)
    input wire [1:0] M_AXI_3_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 ARVALID" *)
    output wire M_AXI_3_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 ARREADY" *)
    input wire M_AXI_3_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 ARADDR" *)
    output wire [32-1:0] M_AXI_3_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 ARPROT" *)
    output wire [2:0] M_AXI_3_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 RVALID" *)
    input wire M_AXI_3_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 RREADY" *)
    output wire M_AXI_3_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 RRESP" *)
    input wire [1:0] M_AXI_3_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_3 RDATA" *)
    input wire [32-1:0] M_AXI_3_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 AWVALID" *)
    output wire M_AXI_4_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 AWREADY" *)
    input wire M_AXI_4_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 AWADDR" *)
    output wire [32-1:0] M_AXI_4_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 AWPROT" *)
    output wire [2:0] M_AXI_4_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 WVALID" *)
    output wire M_AXI_4_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 WREADY" *)
    input wire M_AXI_4_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 WDATA" *)
    output wire [32-1:0] M_AXI_4_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 WSTRB" *)
    output wire [4-1:0] M_AXI_4_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 BVALID" *)
    input wire M_AXI_4_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 BREADY" *)
    output wire M_AXI_4_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 BRESP" *)
    input wire [1:0] M_AXI_4_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 ARVALID" *)
    output wire M_AXI_4_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 ARREADY" *)
    input wire M_AXI_4_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 ARADDR" *)
    output wire [32-1:0] M_AXI_4_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 ARPROT" *)
    output wire [2:0] M_AXI_4_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 RVALID" *)
    input wire M_AXI_4_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 RREADY" *)
    output wire M_AXI_4_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 RRESP" *)
    input wire [1:0] M_AXI_4_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_4 RDATA" *)
    input wire [32-1:0] M_AXI_4_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 AWVALID" *)
    output wire M_AXI_5_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 AWREADY" *)
    input wire M_AXI_5_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 AWADDR" *)
    output wire [32-1:0] M_AXI_5_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 AWPROT" *)
    output wire [2:0] M_AXI_5_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 WVALID" *)
    output wire M_AXI_5_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 WREADY" *)
    input wire M_AXI_5_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 WDATA" *)
    output wire [32-1:0] M_AXI_5_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 WSTRB" *)
    output wire [4-1:0] M_AXI_5_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 BVALID" *)
    input wire M_AXI_5_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 BREADY" *)
    output wire M_AXI_5_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 BRESP" *)
    input wire [1:0] M_AXI_5_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 ARVALID" *)
    output wire M_AXI_5_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 ARREADY" *)
    input wire M_AXI_5_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 ARADDR" *)
    output wire [32-1:0] M_AXI_5_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 ARPROT" *)
    output wire [2:0] M_AXI_5_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 RVALID" *)
    input wire M_AXI_5_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 RREADY" *)
    output wire M_AXI_5_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 RRESP" *)
    input wire [1:0] M_AXI_5_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_5 RDATA" *)
    input wire [32-1:0] M_AXI_5_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 AWVALID" *)
    output wire M_AXI_6_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 AWREADY" *)
    input wire M_AXI_6_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 AWADDR" *)
    output wire [32-1:0] M_AXI_6_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 AWPROT" *)
    output wire [2:0] M_AXI_6_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 WVALID" *)
    output wire M_AXI_6_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 WREADY" *)
    input wire M_AXI_6_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 WDATA" *)
    output wire [32-1:0] M_AXI_6_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 WSTRB" *)
    output wire [4-1:0] M_AXI_6_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 BVALID" *)
    input wire M_AXI_6_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 BREADY" *)
    output wire M_AXI_6_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 BRESP" *)
    input wire [1:0] M_AXI_6_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 ARVALID" *)
    output wire M_AXI_6_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 ARREADY" *)
    input wire M_AXI_6_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 ARADDR" *)
    output wire [32-1:0] M_AXI_6_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 ARPROT" *)
    output wire [2:0] M_AXI_6_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 RVALID" *)
    input wire M_AXI_6_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 RREADY" *)
    output wire M_AXI_6_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 RRESP" *)
    input wire [1:0] M_AXI_6_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_6 RDATA" *)
    input wire [32-1:0] M_AXI_6_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 AWVALID" *)
    output wire M_AXI_7_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 AWREADY" *)
    input wire M_AXI_7_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 AWADDR" *)
    output wire [32-1:0] M_AXI_7_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 AWPROT" *)
    output wire [2:0] M_AXI_7_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 WVALID" *)
    output wire M_AXI_7_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 WREADY" *)
    input wire M_AXI_7_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 WDATA" *)
    output wire [32-1:0] M_AXI_7_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 WSTRB" *)
    output wire [4-1:0] M_AXI_7_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 BVALID" *)
    input wire M_AXI_7_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 BREADY" *)
    output wire M_AXI_7_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 BRESP" *)
    input wire [1:0] M_AXI_7_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 ARVALID" *)
    output wire M_AXI_7_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 ARREADY" *)
    input wire M_AXI_7_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 ARADDR" *)
    output wire [32-1:0] M_AXI_7_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 ARPROT" *)
    output wire [2:0] M_AXI_7_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 RVALID" *)
    input wire M_AXI_7_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 RREADY" *)
    output wire M_AXI_7_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 RRESP" *)
    input wire [1:0] M_AXI_7_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_7 RDATA" *)
    input wire [32-1:0] M_AXI_7_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 AWVALID" *)
    output wire M_AXI_8_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 AWREADY" *)
    input wire M_AXI_8_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 AWADDR" *)
    output wire [32-1:0] M_AXI_8_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 AWPROT" *)
    output wire [2:0] M_AXI_8_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 WVALID" *)
    output wire M_AXI_8_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 WREADY" *)
    input wire M_AXI_8_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 WDATA" *)
    output wire [32-1:0] M_AXI_8_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 WSTRB" *)
    output wire [4-1:0] M_AXI_8_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 BVALID" *)
    input wire M_AXI_8_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 BREADY" *)
    output wire M_AXI_8_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 BRESP" *)
    input wire [1:0] M_AXI_8_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 ARVALID" *)
    output wire M_AXI_8_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 ARREADY" *)
    input wire M_AXI_8_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 ARADDR" *)
    output wire [32-1:0] M_AXI_8_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 ARPROT" *)
    output wire [2:0] M_AXI_8_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 RVALID" *)
    input wire M_AXI_8_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 RREADY" *)
    output wire M_AXI_8_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 RRESP" *)
    input wire [1:0] M_AXI_8_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_8 RDATA" *)
    input wire [32-1:0] M_AXI_8_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 AWVALID" *)
    output wire M_AXI_9_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 AWREADY" *)
    input wire M_AXI_9_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 AWADDR" *)
    output wire [32-1:0] M_AXI_9_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 AWPROT" *)
    output wire [2:0] M_AXI_9_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 WVALID" *)
    output wire M_AXI_9_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 WREADY" *)
    input wire M_AXI_9_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 WDATA" *)
    output wire [32-1:0] M_AXI_9_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 WSTRB" *)
    output wire [4-1:0] M_AXI_9_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 BVALID" *)
    input wire M_AXI_9_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 BREADY" *)
    output wire M_AXI_9_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 BRESP" *)
    input wire [1:0] M_AXI_9_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 ARVALID" *)
    output wire M_AXI_9_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 ARREADY" *)
    input wire M_AXI_9_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 ARADDR" *)
    output wire [32-1:0] M_AXI_9_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 ARPROT" *)
    output wire [2:0] M_AXI_9_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 RVALID" *)
    input wire M_AXI_9_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 RREADY" *)
    output wire M_AXI_9_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 RRESP" *)
    input wire [1:0] M_AXI_9_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_9 RDATA" *)
    input wire [32-1:0] M_AXI_9_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 AWVALID" *)
    output wire M_AXI_10_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 AWREADY" *)
    input wire M_AXI_10_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 AWADDR" *)
    output wire [32-1:0] M_AXI_10_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 AWPROT" *)
    output wire [2:0] M_AXI_10_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 WVALID" *)
    output wire M_AXI_10_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 WREADY" *)
    input wire M_AXI_10_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 WDATA" *)
    output wire [32-1:0] M_AXI_10_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 WSTRB" *)
    output wire [4-1:0] M_AXI_10_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 BVALID" *)
    input wire M_AXI_10_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 BREADY" *)
    output wire M_AXI_10_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 BRESP" *)
    input wire [1:0] M_AXI_10_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 ARVALID" *)
    output wire M_AXI_10_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 ARREADY" *)
    input wire M_AXI_10_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 ARADDR" *)
    output wire [32-1:0] M_AXI_10_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 ARPROT" *)
    output wire [2:0] M_AXI_10_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 RVALID" *)
    input wire M_AXI_10_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 RREADY" *)
    output wire M_AXI_10_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 RRESP" *)
    input wire [1:0] M_AXI_10_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_10 RDATA" *)
    input wire [32-1:0] M_AXI_10_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 AWVALID" *)
    output wire M_AXI_11_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 AWREADY" *)
    input wire M_AXI_11_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 AWADDR" *)
    output wire [32-1:0] M_AXI_11_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 AWPROT" *)
    output wire [2:0] M_AXI_11_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 WVALID" *)
    output wire M_AXI_11_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 WREADY" *)
    input wire M_AXI_11_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 WDATA" *)
    output wire [32-1:0] M_AXI_11_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 WSTRB" *)
    output wire [4-1:0] M_AXI_11_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 BVALID" *)
    input wire M_AXI_11_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 BREADY" *)
    output wire M_AXI_11_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 BRESP" *)
    input wire [1:0] M_AXI_11_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 ARVALID" *)
    output wire M_AXI_11_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 ARREADY" *)
    input wire M_AXI_11_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 ARADDR" *)
    output wire [32-1:0] M_AXI_11_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 ARPROT" *)
    output wire [2:0] M_AXI_11_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 RVALID" *)
    input wire M_AXI_11_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 RREADY" *)
    output wire M_AXI_11_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 RRESP" *)
    input wire [1:0] M_AXI_11_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_11 RDATA" *)
    input wire [32-1:0] M_AXI_11_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 AWVALID" *)
    output wire M_AXI_12_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 AWREADY" *)
    input wire M_AXI_12_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 AWADDR" *)
    output wire [32-1:0] M_AXI_12_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 AWPROT" *)
    output wire [2:0] M_AXI_12_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 WVALID" *)
    output wire M_AXI_12_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 WREADY" *)
    input wire M_AXI_12_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 WDATA" *)
    output wire [32-1:0] M_AXI_12_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 WSTRB" *)
    output wire [4-1:0] M_AXI_12_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 BVALID" *)
    input wire M_AXI_12_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 BREADY" *)
    output wire M_AXI_12_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 BRESP" *)
    input wire [1:0] M_AXI_12_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 ARVALID" *)
    output wire M_AXI_12_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 ARREADY" *)
    input wire M_AXI_12_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 ARADDR" *)
    output wire [32-1:0] M_AXI_12_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 ARPROT" *)
    output wire [2:0] M_AXI_12_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 RVALID" *)
    input wire M_AXI_12_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 RREADY" *)
    output wire M_AXI_12_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 RRESP" *)
    input wire [1:0] M_AXI_12_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_12 RDATA" *)
    input wire [32-1:0] M_AXI_12_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 AWVALID" *)
    output wire M_AXI_13_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 AWREADY" *)
    input wire M_AXI_13_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 AWADDR" *)
    output wire [32-1:0] M_AXI_13_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 AWPROT" *)
    output wire [2:0] M_AXI_13_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 WVALID" *)
    output wire M_AXI_13_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 WREADY" *)
    input wire M_AXI_13_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 WDATA" *)
    output wire [32-1:0] M_AXI_13_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 WSTRB" *)
    output wire [4-1:0] M_AXI_13_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 BVALID" *)
    input wire M_AXI_13_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 BREADY" *)
    output wire M_AXI_13_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 BRESP" *)
    input wire [1:0] M_AXI_13_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 ARVALID" *)
    output wire M_AXI_13_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 ARREADY" *)
    input wire M_AXI_13_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 ARADDR" *)
    output wire [32-1:0] M_AXI_13_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 ARPROT" *)
    output wire [2:0] M_AXI_13_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 RVALID" *)
    input wire M_AXI_13_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 RREADY" *)
    output wire M_AXI_13_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 RRESP" *)
    input wire [1:0] M_AXI_13_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_13 RDATA" *)
    input wire [32-1:0] M_AXI_13_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 AWVALID" *)
    output wire M_AXI_14_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 AWREADY" *)
    input wire M_AXI_14_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 AWADDR" *)
    output wire [32-1:0] M_AXI_14_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 AWPROT" *)
    output wire [2:0] M_AXI_14_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 WVALID" *)
    output wire M_AXI_14_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 WREADY" *)
    input wire M_AXI_14_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 WDATA" *)
    output wire [32-1:0] M_AXI_14_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 WSTRB" *)
    output wire [4-1:0] M_AXI_14_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 BVALID" *)
    input wire M_AXI_14_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 BREADY" *)
    output wire M_AXI_14_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 BRESP" *)
    input wire [1:0] M_AXI_14_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 ARVALID" *)
    output wire M_AXI_14_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 ARREADY" *)
    input wire M_AXI_14_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 ARADDR" *)
    output wire [32-1:0] M_AXI_14_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 ARPROT" *)
    output wire [2:0] M_AXI_14_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 RVALID" *)
    input wire M_AXI_14_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 RREADY" *)
    output wire M_AXI_14_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 RRESP" *)
    input wire [1:0] M_AXI_14_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_14 RDATA" *)
    input wire [32-1:0] M_AXI_14_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 AWVALID" *)
    output wire M_AXI_15_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 AWREADY" *)
    input wire M_AXI_15_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 AWADDR" *)
    output wire [32-1:0] M_AXI_15_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 AWPROT" *)
    output wire [2:0] M_AXI_15_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 WVALID" *)
    output wire M_AXI_15_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 WREADY" *)
    input wire M_AXI_15_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 WDATA" *)
    output wire [32-1:0] M_AXI_15_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 WSTRB" *)
    output wire [4-1:0] M_AXI_15_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 BVALID" *)
    input wire M_AXI_15_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 BREADY" *)
    output wire M_AXI_15_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 BRESP" *)
    input wire [1:0] M_AXI_15_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 ARVALID" *)
    output wire M_AXI_15_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 ARREADY" *)
    input wire M_AXI_15_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 ARADDR" *)
    output wire [32-1:0] M_AXI_15_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 ARPROT" *)
    output wire [2:0] M_AXI_15_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 RVALID" *)
    input wire M_AXI_15_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 RREADY" *)
    output wire M_AXI_15_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 RRESP" *)
    input wire [1:0] M_AXI_15_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 m_axi_15 RDATA" *)
    input wire [32-1:0] M_AXI_15_RDATA,
    
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 AWVALID" *)
    input wire S_AXI_0_AWVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 AWREADY" *)
    output wire S_AXI_0_AWREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 AWADDR" *)
    input wire [32-1:0] S_AXI_0_AWADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 AWPROT" *)
    input wire [2:0] S_AXI_0_AWPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 WVALID" *)
    input wire S_AXI_0_WVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 WREADY" *)
    output wire S_AXI_0_WREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 WDATA" *)
    input wire [32-1:0] S_AXI_0_WDATA,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 WSTRB" *)
    input wire [4-1:0] S_AXI_0_WSTRB,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 BVALID" *)
    output wire S_AXI_0_BVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 BREADY" *)
    input wire S_AXI_0_BREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 BRESP" *)
    output wire [1:0] S_AXI_0_BRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 ARVALID" *)
    input wire S_AXI_0_ARVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 ARREADY" *)
    output wire S_AXI_0_ARREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 ARADDR" *)
    input wire [32-1:0] S_AXI_0_ARADDR,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 ARPROT" *)
    input wire [2:0] S_AXI_0_ARPROT,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 RVALID" *)
    output wire S_AXI_0_RVALID,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 RREADY" *)
    input wire S_AXI_0_RREADY,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 RRESP" *)
    output wire [1:0] S_AXI_0_RRESP,
    (* X_INTERFACE_INFO = "xilinx.com:interface:aximm:1.0 s_axi_0 RDATA" *)
    output wire [32-1:0] S_AXI_0_RDATA
    );
    axilxbar #(
    .C_AXI_DATA_WIDTH(32),
    .C_AXI_ADDR_WIDTH(32),
    .NM(1),
    .NS(16),
    .SLAVE_ADDR(
{32'h0031_0000,
32'h0030_0000,
32'h0022_0000,
32'h0020_0000,
32'h001A_0000,
32'h0019_0000,
32'h0018_0000,
32'h0017_0000,
32'h0016_0000,
32'h0015_0000,
32'h0014_0000,
32'h0013_0000,
32'h0011_0000,
32'h0010_0000,
32'h0002_0000,
32'h0001_0000} ),
    .SLAVE_MASK({16{ 32'h00FF0000 }})
    ) axilxbar_inst (
    .S_AXI_AWVALID({S_AXI_0_AWVALID}),
.S_AXI_AWREADY({S_AXI_0_AWREADY}),
.S_AXI_AWADDR({S_AXI_0_AWADDR}),
.S_AXI_AWPROT({S_AXI_0_AWPROT}),
.S_AXI_WVALID({S_AXI_0_WVALID}),
.S_AXI_WREADY({S_AXI_0_WREADY}),
.S_AXI_WDATA({S_AXI_0_WDATA}),
.S_AXI_WSTRB({S_AXI_0_WSTRB}),
.S_AXI_BVALID({S_AXI_0_BVALID}),
.S_AXI_BREADY({S_AXI_0_BREADY}),
.S_AXI_BRESP({S_AXI_0_BRESP}),
.S_AXI_ARVALID({S_AXI_0_ARVALID}),
.S_AXI_ARREADY({S_AXI_0_ARREADY}),
.S_AXI_ARADDR({S_AXI_0_ARADDR}),
.S_AXI_ARPROT({S_AXI_0_ARPROT}),
.S_AXI_RVALID({S_AXI_0_RVALID}),
.S_AXI_RREADY({S_AXI_0_RREADY}),
.S_AXI_RDATA({S_AXI_0_RDATA}),
.S_AXI_RRESP({S_AXI_0_RRESP}),
.M_AXI_AWVALID({M_AXI_15_AWVALID,M_AXI_14_AWVALID,M_AXI_13_AWVALID,M_AXI_12_AWVALID,M_AXI_11_AWVALID,M_AXI_10_AWVALID,M_AXI_9_AWVALID,M_AXI_8_AWVALID,M_AXI_7_AWVALID,M_AXI_6_AWVALID,M_AXI_5_AWVALID,M_AXI_4_AWVALID,M_AXI_3_AWVALID,M_AXI_2_AWVALID,M_AXI_1_AWVALID,M_AXI_0_AWVALID}),
.M_AXI_AWREADY({M_AXI_15_AWREADY,M_AXI_14_AWREADY,M_AXI_13_AWREADY,M_AXI_12_AWREADY,M_AXI_11_AWREADY,M_AXI_10_AWREADY,M_AXI_9_AWREADY,M_AXI_8_AWREADY,M_AXI_7_AWREADY,M_AXI_6_AWREADY,M_AXI_5_AWREADY,M_AXI_4_AWREADY,M_AXI_3_AWREADY,M_AXI_2_AWREADY,M_AXI_1_AWREADY,M_AXI_0_AWREADY}),
.M_AXI_AWADDR({M_AXI_15_AWADDR,M_AXI_14_AWADDR,M_AXI_13_AWADDR,M_AXI_12_AWADDR,M_AXI_11_AWADDR,M_AXI_10_AWADDR,M_AXI_9_AWADDR,M_AXI_8_AWADDR,M_AXI_7_AWADDR,M_AXI_6_AWADDR,M_AXI_5_AWADDR,M_AXI_4_AWADDR,M_AXI_3_AWADDR,M_AXI_2_AWADDR,M_AXI_1_AWADDR,M_AXI_0_AWADDR}),
.M_AXI_AWPROT({M_AXI_15_AWPROT,M_AXI_14_AWPROT,M_AXI_13_AWPROT,M_AXI_12_AWPROT,M_AXI_11_AWPROT,M_AXI_10_AWPROT,M_AXI_9_AWPROT,M_AXI_8_AWPROT,M_AXI_7_AWPROT,M_AXI_6_AWPROT,M_AXI_5_AWPROT,M_AXI_4_AWPROT,M_AXI_3_AWPROT,M_AXI_2_AWPROT,M_AXI_1_AWPROT,M_AXI_0_AWPROT}),
.M_AXI_WVALID({M_AXI_15_WVALID,M_AXI_14_WVALID,M_AXI_13_WVALID,M_AXI_12_WVALID,M_AXI_11_WVALID,M_AXI_10_WVALID,M_AXI_9_WVALID,M_AXI_8_WVALID,M_AXI_7_WVALID,M_AXI_6_WVALID,M_AXI_5_WVALID,M_AXI_4_WVALID,M_AXI_3_WVALID,M_AXI_2_WVALID,M_AXI_1_WVALID,M_AXI_0_WVALID}),
.M_AXI_WREADY({M_AXI_15_WREADY,M_AXI_14_WREADY,M_AXI_13_WREADY,M_AXI_12_WREADY,M_AXI_11_WREADY,M_AXI_10_WREADY,M_AXI_9_WREADY,M_AXI_8_WREADY,M_AXI_7_WREADY,M_AXI_6_WREADY,M_AXI_5_WREADY,M_AXI_4_WREADY,M_AXI_3_WREADY,M_AXI_2_WREADY,M_AXI_1_WREADY,M_AXI_0_WREADY}),
.M_AXI_WDATA({M_AXI_15_WDATA,M_AXI_14_WDATA,M_AXI_13_WDATA,M_AXI_12_WDATA,M_AXI_11_WDATA,M_AXI_10_WDATA,M_AXI_9_WDATA,M_AXI_8_WDATA,M_AXI_7_WDATA,M_AXI_6_WDATA,M_AXI_5_WDATA,M_AXI_4_WDATA,M_AXI_3_WDATA,M_AXI_2_WDATA,M_AXI_1_WDATA,M_AXI_0_WDATA}),
.M_AXI_WSTRB({M_AXI_15_WSTRB,M_AXI_14_WSTRB,M_AXI_13_WSTRB,M_AXI_12_WSTRB,M_AXI_11_WSTRB,M_AXI_10_WSTRB,M_AXI_9_WSTRB,M_AXI_8_WSTRB,M_AXI_7_WSTRB,M_AXI_6_WSTRB,M_AXI_5_WSTRB,M_AXI_4_WSTRB,M_AXI_3_WSTRB,M_AXI_2_WSTRB,M_AXI_1_WSTRB,M_AXI_0_WSTRB}),
.M_AXI_BVALID({M_AXI_15_BVALID,M_AXI_14_BVALID,M_AXI_13_BVALID,M_AXI_12_BVALID,M_AXI_11_BVALID,M_AXI_10_BVALID,M_AXI_9_BVALID,M_AXI_8_BVALID,M_AXI_7_BVALID,M_AXI_6_BVALID,M_AXI_5_BVALID,M_AXI_4_BVALID,M_AXI_3_BVALID,M_AXI_2_BVALID,M_AXI_1_BVALID,M_AXI_0_BVALID}),
.M_AXI_BREADY({M_AXI_15_BREADY,M_AXI_14_BREADY,M_AXI_13_BREADY,M_AXI_12_BREADY,M_AXI_11_BREADY,M_AXI_10_BREADY,M_AXI_9_BREADY,M_AXI_8_BREADY,M_AXI_7_BREADY,M_AXI_6_BREADY,M_AXI_5_BREADY,M_AXI_4_BREADY,M_AXI_3_BREADY,M_AXI_2_BREADY,M_AXI_1_BREADY,M_AXI_0_BREADY}),
.M_AXI_BRESP({M_AXI_15_BRESP,M_AXI_14_BRESP,M_AXI_13_BRESP,M_AXI_12_BRESP,M_AXI_11_BRESP,M_AXI_10_BRESP,M_AXI_9_BRESP,M_AXI_8_BRESP,M_AXI_7_BRESP,M_AXI_6_BRESP,M_AXI_5_BRESP,M_AXI_4_BRESP,M_AXI_3_BRESP,M_AXI_2_BRESP,M_AXI_1_BRESP,M_AXI_0_BRESP}),
.M_AXI_ARVALID({M_AXI_15_ARVALID,M_AXI_14_ARVALID,M_AXI_13_ARVALID,M_AXI_12_ARVALID,M_AXI_11_ARVALID,M_AXI_10_ARVALID,M_AXI_9_ARVALID,M_AXI_8_ARVALID,M_AXI_7_ARVALID,M_AXI_6_ARVALID,M_AXI_5_ARVALID,M_AXI_4_ARVALID,M_AXI_3_ARVALID,M_AXI_2_ARVALID,M_AXI_1_ARVALID,M_AXI_0_ARVALID}),
.M_AXI_ARREADY({M_AXI_15_ARREADY,M_AXI_14_ARREADY,M_AXI_13_ARREADY,M_AXI_12_ARREADY,M_AXI_11_ARREADY,M_AXI_10_ARREADY,M_AXI_9_ARREADY,M_AXI_8_ARREADY,M_AXI_7_ARREADY,M_AXI_6_ARREADY,M_AXI_5_ARREADY,M_AXI_4_ARREADY,M_AXI_3_ARREADY,M_AXI_2_ARREADY,M_AXI_1_ARREADY,M_AXI_0_ARREADY}),
.M_AXI_ARADDR({M_AXI_15_ARADDR,M_AXI_14_ARADDR,M_AXI_13_ARADDR,M_AXI_12_ARADDR,M_AXI_11_ARADDR,M_AXI_10_ARADDR,M_AXI_9_ARADDR,M_AXI_8_ARADDR,M_AXI_7_ARADDR,M_AXI_6_ARADDR,M_AXI_5_ARADDR,M_AXI_4_ARADDR,M_AXI_3_ARADDR,M_AXI_2_ARADDR,M_AXI_1_ARADDR,M_AXI_0_ARADDR}),
.M_AXI_ARPROT({M_AXI_15_ARPROT,M_AXI_14_ARPROT,M_AXI_13_ARPROT,M_AXI_12_ARPROT,M_AXI_11_ARPROT,M_AXI_10_ARPROT,M_AXI_9_ARPROT,M_AXI_8_ARPROT,M_AXI_7_ARPROT,M_AXI_6_ARPROT,M_AXI_5_ARPROT,M_AXI_4_ARPROT,M_AXI_3_ARPROT,M_AXI_2_ARPROT,M_AXI_1_ARPROT,M_AXI_0_ARPROT}),
.M_AXI_RVALID({M_AXI_15_RVALID,M_AXI_14_RVALID,M_AXI_13_RVALID,M_AXI_12_RVALID,M_AXI_11_RVALID,M_AXI_10_RVALID,M_AXI_9_RVALID,M_AXI_8_RVALID,M_AXI_7_RVALID,M_AXI_6_RVALID,M_AXI_5_RVALID,M_AXI_4_RVALID,M_AXI_3_RVALID,M_AXI_2_RVALID,M_AXI_1_RVALID,M_AXI_0_RVALID}),
.M_AXI_RREADY({M_AXI_15_RREADY,M_AXI_14_RREADY,M_AXI_13_RREADY,M_AXI_12_RREADY,M_AXI_11_RREADY,M_AXI_10_RREADY,M_AXI_9_RREADY,M_AXI_8_RREADY,M_AXI_7_RREADY,M_AXI_6_RREADY,M_AXI_5_RREADY,M_AXI_4_RREADY,M_AXI_3_RREADY,M_AXI_2_RREADY,M_AXI_1_RREADY,M_AXI_0_RREADY}),
.M_AXI_RDATA({M_AXI_15_RDATA,M_AXI_14_RDATA,M_AXI_13_RDATA,M_AXI_12_RDATA,M_AXI_11_RDATA,M_AXI_10_RDATA,M_AXI_9_RDATA,M_AXI_8_RDATA,M_AXI_7_RDATA,M_AXI_6_RDATA,M_AXI_5_RDATA,M_AXI_4_RDATA,M_AXI_3_RDATA,M_AXI_2_RDATA,M_AXI_1_RDATA,M_AXI_0_RDATA}),
.M_AXI_RRESP({M_AXI_15_RRESP,M_AXI_14_RRESP,M_AXI_13_RRESP,M_AXI_12_RRESP,M_AXI_11_RRESP,M_AXI_10_RRESP,M_AXI_9_RRESP,M_AXI_8_RRESP,M_AXI_7_RRESP,M_AXI_6_RRESP,M_AXI_5_RRESP,M_AXI_4_RRESP,M_AXI_3_RRESP,M_AXI_2_RRESP,M_AXI_1_RRESP,M_AXI_0_RRESP}),

    .S_AXI_ACLK(S_AXI_ACLK),
    .S_AXI_ARESETN(S_AXI_ARESETN)
    );
    endmodule
    